 LIBRARY IEEE ;
 USE IEEE.STD_LOGIC_1164.ALL ;
 ENTITY DECL7S IS
  PORT ( A  : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
      LED7S : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)  ) ;
 END ;
 ARCHITECTURE one OF DECL7S IS
 BEGIN
  PROCESS( A )
  BEGIN
  CASE  A  IS
   WHEN "0000" =>  LED7S <= "0111111" ; 
   WHEN "0001" =>  LED7S <= "0000110" ; 
   WHEN "0010" =>  LED7S <= "1011011" ; 
   WHEN "0011" =>  LED7S <= "1001111" ; 
   WHEN "0100" =>  LED7S <= "1100110" ; 
   WHEN "0101" =>  LED7S <= "1101101" ; 
   WHEN "0110" =>  LED7S <= "1111101" ;
   WHEN "0111" =>  LED7S <= "0000111" ;
   WHEN "1000" =>  LED7S <= "1111111" ; 
   WHEN "1001" =>  LED7S <= "1101111" ; 
   WHEN "1010" =>  LED7S <= "1110111" ; 
   WHEN "1011" =>  LED7S <= "1111100" ;
   WHEN "1100" =>  LED7S <= "0111001" ;
   WHEN "1101" =>  LED7S <= "1011110" ; 
   WHEN "1110" =>  LED7S <= "1111001" ;
   WHEN "1111" =>  LED7S <= "1110001" ;
   WHEN OTHERS =>  NULL ;
   END CASE ;
  END PROCESS ;
 END ;
