library verilog;
use verilog.vl_types.all;
entity step_vlg_vec_tst is
end step_vlg_vec_tst;
