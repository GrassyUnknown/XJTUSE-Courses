library verilog;
use verilog.vl_types.all;
entity step2_vlg_vec_tst is
end step2_vlg_vec_tst;
