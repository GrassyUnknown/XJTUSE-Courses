library verilog;
use verilog.vl_types.all;
entity PC_vlg_vec_tst is
end PC_vlg_vec_tst;
