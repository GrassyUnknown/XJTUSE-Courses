LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY REG8 IS
    PORT (  Load :  IN STD_LOGIC;
             A  :  IN STD_LOGIC_VECTOR(7 DOWNTO 0);
             B  : OUT STD_LOGIC_VECTOR(7 DOWNTO 0) );
END REG8;
ARCHITECTURE behav OF REG8 IS
BEGIN
    PROCESS(Load, A)
   BEGIN
   IF Load'EVENT AND Load = '1' THEN   
            B <= A; 
        END IF;
    END PROCESS;
END behav;


