library verilog;
use verilog.vl_types.all;
entity exp2_2_vlg_vec_tst is
end exp2_2_vlg_vec_tst;
