library verilog;
use verilog.vl_types.all;
entity step3_vlg_vec_tst is
end step3_vlg_vec_tst;
