library verilog;
use verilog.vl_types.all;
entity ALU_vlg_vec_tst is
end ALU_vlg_vec_tst;
