 LIBRARY IEEE ;
 USE IEEE.STD_LOGIC_1164.ALL ;
 ENTITY MUX48 IS
  PORT (   S  : IN  STD_LOGIC_VECTOR(2 DOWNTO 0);
           A1 : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
           A2 : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
           A3 : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
           A4 : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
           A5 : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
           A6 : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
           A7 : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
           A8 : IN  STD_LOGIC_VECTOR(3 DOWNTO 0);
           RT : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)   ) ;
 END ;
 ARCHITECTURE one OF MUX48 IS
 BEGIN
  RT <= A1 WHEN S= "111"  ELSE
        A2 WHEN S= "110"  ELSE
        A3 WHEN S= "101"  ELSE
        A4 WHEN S= "100"  ELSE
        A5 WHEN S= "011"  ELSE
        A6 WHEN S= "010"  ELSE
        A7 WHEN S= "001"  ELSE
        A8 WHEN S= "000"  ELSE
        A8 ;
 END ;
