library verilog;
use verilog.vl_types.all;
entity LDR0_2_vlg_vec_tst is
end LDR0_2_vlg_vec_tst;
