library verilog;
use verilog.vl_types.all;
entity uA_reg_vlg_vec_tst is
end uA_reg_vlg_vec_tst;
