LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY REG10B IS
    PORT (  Load :  IN STD_LOGIC;
             DIN :  IN STD_LOGIC_VECTOR(9 DOWNTO 0);
            DOUT : OUT STD_LOGIC_VECTOR(9 DOWNTO 0) );
END REG10B;
ARCHITECTURE behav OF REG10B IS
BEGIN
    PROCESS(Load, DIN)
   BEGIN
   IF Load'EVENT AND Load = '1' THEN    -- ʱ�ӵ���ʱ��������������
            DOUT <= DIN;
        END IF;
    END PROCESS;
END behav;


