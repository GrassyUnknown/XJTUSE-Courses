library verilog;
use verilog.vl_types.all;
entity AR_vlg_vec_tst is
end AR_vlg_vec_tst;
