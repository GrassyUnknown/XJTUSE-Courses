LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
ENTITY ADDER32B IS
    PORT (  A : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
            B : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
            S : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)     );
END ADDER32B;
ARCHITECTURE behav OF ADDER32B IS
    BEGIN
	S <= A + B;
END behav;


