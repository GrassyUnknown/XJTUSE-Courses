library verilog;
use verilog.vl_types.all;
entity exp2_1_vlg_check_tst is
    port(
        q               : in     vl_logic_vector(23 downto 0);
        sampler_rx      : in     vl_logic
    );
end exp2_1_vlg_check_tst;
